library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity control_memory is
    Port ( 
       CAR_in : in std_logic_vector(7 downto 0);
       NA : out  std_logic_vector(7 downto 0);
       MS : out  std_logic_vector(2 downto 0);
       FS : out std_logic_vector(4 downto 0);
       MC,IL,PI,PL,TD,TA,TB,MB,MD,RW,MM,MW : out std_logic
    );
end control_memory;

architecture Behavioral of control_memory is
type mem_array is array(0 to 255) of std_logic_vector(27 downto 0);

begin
memory_m: process(CAR_in)
variable control_mem : mem_array:=(
    x"C020306", 
    x"C02400E",	
    x"C020184",
    X"0000000",
    X"0000000", 
    X"0000000", 
    X"0000000", 
    X"0000000", 
    X"0000000", 
    X"0000000", 
    X"0000000", 
    X"0000000", 
    --12
    X"C020306",
    X"0000000",
    X"0000000", 
    X"0000000", 

    X"C030024", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000",
    
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 

    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000",

    -- 0x60
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 

    -- 0x70
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000",
    
    -- 0x60
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 

    --0x70
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000",
    
    --0x80
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 

    --0x90
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000",
    
    --0xA0
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 

    --0xB0
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000",

    --0xC0
    x"C12C002", x"0030000", X"0000000", X"0000000",
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000",

    --0xD0
    X"C10C002", X"0030004", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000",
    
    --0xE0
    X"C12C002", X"0030000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 

    --0xF0
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000", 
    X"0000000", X"0000000", X"0000000", X"0000000");

    variable addr : integer;
    variable control_out : std_logic_vector(27 downto 0);
begin
    addr := conv_integer(CAR_in);
    control_out := control_mem(addr);
    MW <= control_out(0);
    MM <= control_out(1);
    RW <= control_out(2);
    MD <= control_out(3);
    FS <= control_out(8 downto 4);
    MB <= control_out(9);
    TB <= control_out(10);
    TA <= control_out(11);
    TD <= control_out(12);
    PL <= control_out(13);
    PI <= control_out(14);
    IL <= control_out(15);
    MC <= control_out(16);
    MS <= control_out(19 downto 17);
    NA <= control_out(27 downto 20);
    end process;
end Behavioral;
